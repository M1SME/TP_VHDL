  --Example instantiation for system 'unnamed'
  unnamed_inst : unnamed
    port map(
      Leds_from_the_Anemometre_0 => Leds_from_the_Anemometre_0,
      out_pwm_from_the_avalon_pwm_0 => out_pwm_from_the_avalon_pwm_0,
      IN_PWM_COMPAS_to_the_Anemometre_0 => IN_PWM_COMPAS_to_the_Anemometre_0,
      clk_0 => clk_0,
      reset_n => reset_n
    );


