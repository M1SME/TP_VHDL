  --Example instantiation for system 'mon_SOPC'
  mon_SOPC_inst : mon_SOPC
    port map(
      out_port_from_the_OutputPIO => out_port_from_the_OutputPIO,
      out_pwm_from_the_avalon_pwm_0 => out_pwm_from_the_avalon_pwm_0,
      clk_0 => clk_0,
      in_port_to_the_InputPIO => in_port_to_the_InputPIO,
      reset_n => reset_n
    );


