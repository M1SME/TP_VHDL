  --Example instantiation for system 'CPU_GestionVerin'
  CPU_GestionVerin_inst : CPU_GestionVerin
    port map(
      clk_adc_from_the_GestionVerin_0 => clk_adc_from_the_GestionVerin_0,
      cs_n_from_the_GestionVerin_0 => cs_n_from_the_GestionVerin_0,
      out_PWM_from_the_GestionVerin_0 => out_PWM_from_the_GestionVerin_0,
      out_sens_from_the_GestionVerin_0 => out_sens_from_the_GestionVerin_0,
      Data_IN_to_the_GestionVerin_0 => Data_IN_to_the_GestionVerin_0,
      clk_0 => clk_0,
      reset_n => reset_n
    );


