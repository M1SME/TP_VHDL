  --Example instantiation for system 'CPU_NMEA'
  CPU_NMEA_inst : CPU_NMEA
    port map(
      LEDs_from_the_NMEA_Interface_0 => LEDs_from_the_NMEA_Interface_0,
      Tx_Pin_from_the_NMEA_Interface_0 => Tx_Pin_from_the_NMEA_Interface_0,
      Rx_Pin_to_the_NMEA_Interface_0 => Rx_Pin_to_the_NMEA_Interface_0,
      clk_0 => clk_0,
      reset_n => reset_n
    );


